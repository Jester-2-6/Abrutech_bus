/*
Module name  : bus_top_module.v
Author 	     : W.M.R.R.Wickramasinghe
Date Modified: 06/06/2019
Organization : ABruTECH
Description  : Top module containig the arbiter,masters and slaves
*/

module bus_top_module(
    rstn,
    clk,
    tx0,
    rx0,
    tx1,
    rx1,
    hex0,
    hex1,
    hex2,
    hex3,
    hex4,
    requests,
    utilization,
    slave_busy,
    mux_switch
);

// Parameters

// Port declaration



endmodule