/*
Module name  : serial_parallel.v
Author 	     : W.M.R.R.Wickramasinghe
Date Modified: 01/06/2019
Organization : ABruTECH
Description  : Master module of the bus
*/

module #()serial_parallel(
    clk,
    rstn,
    din,
    dv_in,
    dout,
    dv_out,
    bit_lngt,
    en
);

endmodule